/*
 * Module Name: constant_addition_layer
 * Author(s):
 * Description:
 * Ref: NIST SP 800-232
 */

import ascon_pkg::*;

module constant_addition_layer (
    input   ascon_state_t   state_array_i,
    output  ascon_state_t   state_array_o
);



endmodule
