`timescale 1ns/1ps
import ascon_pkg::*;

module tb_linear_diffusion_layer;

    // DUT signals
    ascon_state_t state_i;
    ascon_state_t state_o;

    // Reference full 320-bit values
    logic [319:0] input_vec;
    logic [319:0] expected_vec;

    // DUT
    linear_diffusion_layer dut (
        .state_array_i(state_i),
        .state_array_o(state_o)
    );

    initial begin
        $display("=== Linear Diffusion Layer Testbench ===");

        // -------------------------
        // Test Vector 1
        // -------------------------
        input_vec =
            320'b01001100001110111000010001000110111100110101111101000100010000100011010111100100101110101110111011101011101010110011101010100011001011101100100001110011001110011011111011010101010100001111011111101100110110111011111001111111001000100100111110111100011000101100110001111101111100000101101001010110111111111011101110000010;
        expected_vec =
            320'b11101011110110100101110011101100010111111001111111100111000010000000000001111000010110010011001000001101011001101010010110111000011001010001011101101011011010011000011101000100101011011100111101110100010000101101001011111110111101011110101111101000000010010101010011110110000100011111100100101111001010111111010011111000;
        state_i = input_vec;
        #1;

        assert (state_o == expected_vec)
            else $fatal(1, "❌ Test Vector 1 FAILED");

        $display("✅ Test Vector 1 PASSED");

        // -------------------------
        // Test Vector 2
        // -------------------------
        input_vec =
            320'b01111001000000010101111000110110000110111100111010101011000111100010101111101010101110001101010011101100001101000110010001011000111110111010001001010000101110000001100111010110011010000011001000001010000000100001000111110001110011010000000110010100101100000000000110100100110111100010111000010111010000011000000000101101;

        expected_vec =
            320'b01011110111111101011101111011111111110001100010110110110111001110000111111001100010101111000111110000101011001010001111101011011010011011001110111110001101001101111010101011010000001011000101110111001100010001001110101010110110001010001100100110101000100110100010110111001011111001100101010010110110010011010000000100100;
        state_i = input_vec;
        #1;

        assert (state_o == expected_vec)
            else $fatal(1, "❌ Test Vector  FAILED");

        $display("✅ Test Vector 2 PASSED");

        $display("🎉 All tests PASSED");
        $finish;
    end

endmodule
